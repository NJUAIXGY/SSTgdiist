module test;
  initial begin
    $display("Hello, Verilog!");
    $finish;
  end
endmodule